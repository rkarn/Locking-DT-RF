`timescale 1ns / 1ps
//Correct KEY=[1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1]
module decision(
KEY,
	feat_8,
	feat_13,
	feat_10,
	feat_12,
	feat_2,
	feat_14,
	feat_9,
	feat_11,
	feat_17,
	feat_16,
	feat_5,
	feat_0,
	feat_1,
	feat_6,
	feat_7,
	feat_3,
	feat_15,
	CLK,
	RST,
	decision
);


	input [9:0] feat_8;
	input [9:0] feat_13;
	input [9:0] feat_10;
	input [9:0] feat_12;
	input [1:0] feat_2;
	input [9:0] feat_14;
	input [9:0] feat_9;
	input [9:0] feat_11;
	input [9:0] feat_17;
	input [9:0] feat_16;
	input [1:0] feat_5;
	input [1:0] feat_0;
	input wire feat_1;
	input [9:0] feat_6;
	input [9:0] feat_7;
	input [1:0] feat_3;
	input [9:0] feat_15;
	input wire CLK;
	input wire RST;
	output [4:0] decision;
input [170:0] KEY;

	wire [9:0] reg_feat_8;
	wire [9:0] reg_feat_13;
	wire [9:0] reg_feat_10;
	wire [9:0] reg_feat_12;
	wire [1:0] reg_feat_2;
	wire [9:0] reg_feat_14;
	wire [9:0] reg_feat_9;
	wire [9:0] reg_feat_11;
	wire [9:0] reg_feat_17;
	wire [9:0] reg_feat_16;
	wire [1:0] reg_feat_5;
	wire [1:0] reg_feat_0;
	wire [0:0] reg_feat_1;
	wire [9:0] reg_feat_6;
	wire [9:0] reg_feat_7;
	wire [1:0] reg_feat_3;
	wire [9:0] reg_feat_15;
	wire [4:0] reg_decision;

wire [0:0] comp_feat_8_538;
wire [0:0] comp_feat_13_632;
wire [0:0] comp_feat_10_734;
wire [0:0] comp_feat_12_453;
wire [0:0] comp_feat_2_2;
wire [0:0] comp_feat_14_504;
wire [0:0] comp_feat_9_6;
wire [0:0] comp_feat_11_744;
wire [0:0] comp_feat_12_240;
wire [0:0] comp_feat_11_823;
wire [0:0] comp_feat_17_787;
wire [0:0] comp_feat_11_742;
wire [0:0] comp_feat_17_765;
wire [0:0] comp_feat_14_537;
wire [0:0] comp_feat_8_506;
wire [0:0] comp_feat_16_741;
wire [0:0] comp_feat_8_491;
wire [0:0] comp_feat_14_535;
wire [0:0] comp_feat_5_2;
wire [0:0] comp_feat_14_525;
wire [0:0] comp_feat_12_537;
wire [0:0] comp_feat_13_626;
wire [0:0] comp_feat_8_512;
wire [0:0] comp_feat_12_523;
wire [0:0] comp_feat_0_0;
wire [0:0] comp_feat_13_608;
wire [0:0] comp_feat_14_522;
wire [0:0] comp_feat_11_770;
wire [0:0] comp_feat_12_517;
wire [0:0] comp_feat_1_0;
wire [0:0] comp_feat_13_538;
wire [0:0] comp_feat_9_356;
wire [0:0] comp_feat_12_526;
wire [0:0] comp_feat_6_359;
wire [0:0] comp_feat_7_480;
wire [0:0] comp_feat_2_1;
wire [0:0] comp_feat_14_512;
wire [0:0] comp_feat_11_763;
wire [0:0] comp_feat_10_696;
wire [0:0] comp_feat_14_502;
wire [0:0] comp_feat_3_0;
wire [0:0] comp_feat_13_588;
wire [0:0] comp_feat_7_469;
wire [0:0] comp_feat_12_493;
wire [0:0] comp_feat_12_486;
wire [0:0] comp_feat_12_512;
wire [0:0] comp_feat_10_752;
wire [0:0] comp_feat_11_727;
wire [0:0] comp_feat_8_493;
wire [0:0] comp_feat_10_767;
wire [0:0] comp_feat_13_623;
wire [0:0] comp_feat_8_510;
wire [0:0] comp_feat_14_487;
wire [0:0] comp_feat_16_685;
wire [0:0] comp_feat_11_728;
wire [0:0] comp_feat_11_718;
wire [0:0] comp_feat_12_490;
wire [0:0] comp_feat_12_504;
wire [0:0] comp_feat_9_508;
wire [0:0] comp_feat_8_524;
wire [0:0] comp_feat_14_499;
wire [0:0] comp_feat_14_495;
wire [0:0] comp_feat_15_856;
wire [0:0] comp_feat_8_461;
wire [0:0] comp_feat_8_452;
wire [0:0] comp_feat_13_627;
wire [0:0] comp_feat_17_767;
wire [0:0] comp_feat_15_787;
wire [0:0] comp_feat_17_752;
wire [0:0] comp_feat_8_475;
wire [0:0] comp_feat_6_361;
wire [0:0] comp_feat_12_521;
wire [0:0] comp_feat_14_521;
wire [0:0] comp_feat_15_803;
wire [0:0] comp_feat_15_732;
wire [0:0] comp_feat_13_612;
wire [0:0] comp_feat_14_509;
wire [0:0] comp_feat_11_719;
wire [0:0] comp_feat_11_693;
wire [0:0] comp_feat_10_772;
wire [0:0] comp_feat_7_487;
wire [0:0] comp_feat_13_573;
wire [0:0] comp_feat_15_820;
wire [0:0] comp_feat_10_775;
wire [0:0] comp_feat_17_862;
wire [0:0] comp_feat_14_531;
wire [0:0] comp_feat_12_515;
wire [0:0] comp_feat_13_606;
wire [0:0] comp_feat_12_528;
wire [0:0] comp_feat_8_528;
wire [0:0] comp_feat_13_633;
wire [0:0] comp_feat_10_759;
wire [0:0] comp_feat_17_841;
wire [0:0] comp_feat_10_0;
wire [0:0] comp_feat_15_863;
wire [0:0] comp_feat_16_702;
wire [0:0] comp_feat_10_770;
wire [0:0] comp_feat_8_487;
wire [0:0] comp_feat_7_470;
wire [0:0] comp_feat_16_735;
wire [0:0] comp_feat_15_781;
wire [0:0] comp_feat_0_1;
wire [0:0] comp_feat_9_533;
wire [0:0] comp_feat_9_536;
wire [0:0] comp_feat_9_826;
wire [0:0] comp_feat_17_827;
wire [0:0] comp_feat_13_636;
wire [0:0] comp_feat_10_749;
wire [0:0] comp_feat_15_648;
wire [0:0] comp_feat_7_388;
wire [0:0] comp_feat_12_525;
wire [0:0] comp_feat_16_684;
wire [0:0] comp_feat_8_462;
wire [0:0] comp_feat_16_751;
wire [0:0] comp_feat_15_892;
wire [0:0] comp_feat_15_747;
wire [0:0] comp_feat_15_640;
wire [0:0] comp_feat_5_1;
wire [0:0] comp_feat_8_401;
wire [0:0] comp_feat_15_741;
wire [0:0] comp_feat_13_938;
wire [0:0] comp_feat_14_520;
wire [0:0] comp_feat_10_689;
wire [0:0] comp_feat_15_756;
wire [0:0] comp_feat_14_493;
wire [0:0] comp_feat_6_396;
wire [0:0] comp_feat_13_647;
wire [0:0] comp_feat_15_823;
wire [0:0] comp_feat_3_1;
wire [0:0] comp_feat_7_472;
wire [0:0] comp_feat_12_518;
wire [0:0] comp_feat_9_515;
wire [0:0] comp_feat_17_833;
wire [0:0] comp_feat_14_505;
wire [0:0] comp_feat_14_526;
wire [0:0] comp_feat_11_831;
wire [0:0] comp_feat_10_712;
wire [0:0] comp_feat_9_213;
wire [0:0] comp_feat_11_837;
wire [0:0] comp_feat_7_464;
wire [0:0] comp_feat_16_731;
wire [0:0] comp_feat_14_23;
wire [0:0] comp_feat_12_536;
wire [0:0] comp_feat_14_529;
wire [0:0] comp_feat_6_409;
wire [0:0] comp_feat_9_511;
wire [0:0] comp_feat_6_385;
wire [0:0] comp_feat_12_520;
wire [0:0] comp_feat_7_476;
wire [0:0] comp_feat_12_497;
wire [0:0] comp_feat_10_755;
wire [0:0] comp_feat_13_614;
wire [0:0] comp_feat_6_378;
wire [0:0] comp_feat_13_582;
wire [0:0] comp_feat_17_763;
wire [0:0] comp_feat_13_628;
wire [0:0] comp_feat_14_566;
wire [0:0] comp_feat_14_536;
wire [0:0] comp_feat_11_827;
wire [0:0] comp_feat_9_558;
wire [0:0] comp_feat_12_533;
wire [0:0] comp_feat_13_613;
wire [0:0] comp_feat_13_574;
wire [0:0] comp_feat_11_753;
wire [0:0] comp_feat_8_542;
wire [0:0] comp_feat_10_753;
wire [0:0] comp_feat_15_806;
wire [0:0] comp_feat_10_676;
wire [0:0] comp_feat_11_410;
wire [0:0] comp_feat_8_586;
wire [0:0] comp_feat_12_431;
COMPS INST_COMP(
KEY,
reg_feat_8, reg_feat_13, reg_feat_10, reg_feat_12, reg_feat_2, reg_feat_14, reg_feat_9, reg_feat_11, reg_feat_17, reg_feat_16, reg_feat_5, reg_feat_0, reg_feat_1, reg_feat_6, reg_feat_7, reg_feat_3, reg_feat_15, comp_feat_8_538, comp_feat_13_632, comp_feat_10_734, comp_feat_12_453, comp_feat_2_2, comp_feat_14_504, comp_feat_9_6, comp_feat_11_744, comp_feat_12_240, comp_feat_11_823, comp_feat_17_787, comp_feat_11_742, comp_feat_17_765, comp_feat_14_537, comp_feat_8_506, comp_feat_16_741, comp_feat_8_491, comp_feat_14_535, comp_feat_5_2, comp_feat_14_525, comp_feat_12_537, comp_feat_13_626, comp_feat_8_512, comp_feat_12_523, comp_feat_0_0, comp_feat_13_608, comp_feat_14_522, comp_feat_11_770, comp_feat_12_517, comp_feat_1_0, comp_feat_13_538, comp_feat_9_356, comp_feat_12_526, comp_feat_6_359, comp_feat_7_480, comp_feat_2_1, comp_feat_14_512, comp_feat_11_763, comp_feat_10_696, comp_feat_14_502, comp_feat_3_0, comp_feat_13_588, comp_feat_7_469, comp_feat_12_493, comp_feat_12_486, comp_feat_12_512, comp_feat_10_752, comp_feat_11_727, comp_feat_8_493, comp_feat_10_767, comp_feat_13_623, comp_feat_8_510, comp_feat_14_487, comp_feat_16_685, comp_feat_11_728, comp_feat_11_718, comp_feat_12_490, comp_feat_12_504, comp_feat_9_508, comp_feat_8_524, comp_feat_14_499, comp_feat_14_495, comp_feat_15_856, comp_feat_8_461, comp_feat_8_452, comp_feat_13_627, comp_feat_17_767, comp_feat_15_787, comp_feat_17_752, comp_feat_8_475, comp_feat_6_361, comp_feat_12_521, comp_feat_14_521, comp_feat_15_803, comp_feat_15_732, comp_feat_13_612, comp_feat_14_509, comp_feat_11_719, comp_feat_11_693, comp_feat_10_772, comp_feat_7_487, comp_feat_13_573, comp_feat_15_820, comp_feat_10_775, comp_feat_17_862, comp_feat_14_531, comp_feat_12_515, comp_feat_13_606, comp_feat_12_528, comp_feat_8_528, comp_feat_13_633, comp_feat_10_759, comp_feat_17_841, comp_feat_10_0, comp_feat_15_863, comp_feat_16_702, comp_feat_10_770, comp_feat_8_487, comp_feat_7_470, comp_feat_16_735, comp_feat_15_781, comp_feat_0_1, comp_feat_9_533, comp_feat_9_536, comp_feat_9_826, comp_feat_17_827, comp_feat_13_636, comp_feat_10_749, comp_feat_15_648, comp_feat_7_388, comp_feat_12_525, comp_feat_16_684, comp_feat_8_462, comp_feat_16_751, comp_feat_15_892, comp_feat_15_747, comp_feat_15_640, comp_feat_5_1, comp_feat_8_401, comp_feat_15_741, comp_feat_13_938, comp_feat_14_520, comp_feat_10_689, comp_feat_15_756, comp_feat_14_493, comp_feat_6_396, comp_feat_13_647, comp_feat_15_823, comp_feat_3_1, comp_feat_7_472, comp_feat_12_518, comp_feat_9_515, comp_feat_17_833, comp_feat_14_505, comp_feat_14_526, comp_feat_11_831, comp_feat_10_712, comp_feat_9_213, comp_feat_11_837, comp_feat_7_464, comp_feat_16_731, comp_feat_14_23, comp_feat_12_536, comp_feat_14_529, comp_feat_6_409, comp_feat_9_511, comp_feat_6_385, comp_feat_12_520, comp_feat_7_476, comp_feat_12_497, comp_feat_10_755, comp_feat_13_614, comp_feat_6_378, comp_feat_13_582, comp_feat_17_763, comp_feat_13_628, comp_feat_14_566, comp_feat_14_536, comp_feat_11_827, comp_feat_9_558, comp_feat_12_533, comp_feat_13_613, comp_feat_13_574, comp_feat_11_753, comp_feat_8_542, comp_feat_10_753, comp_feat_15_806, comp_feat_10_676, comp_feat_11_410, comp_feat_8_586, comp_feat_12_431
);

ANDS INST_ANDS(
comp_feat_8_538, comp_feat_13_632, comp_feat_10_734, comp_feat_12_453, comp_feat_2_2, comp_feat_14_504, comp_feat_9_6, comp_feat_11_744, comp_feat_12_240, comp_feat_11_823, comp_feat_17_787, comp_feat_11_742, comp_feat_17_765, comp_feat_14_537, comp_feat_8_506, comp_feat_16_741, comp_feat_8_491, comp_feat_14_535, comp_feat_5_2, comp_feat_14_525, comp_feat_12_537, comp_feat_13_626, comp_feat_8_512, comp_feat_12_523, comp_feat_0_0, comp_feat_13_608, comp_feat_14_522, comp_feat_11_770, comp_feat_12_517, comp_feat_1_0, comp_feat_13_538, comp_feat_9_356, comp_feat_12_526, comp_feat_6_359, comp_feat_7_480, comp_feat_2_1, comp_feat_14_512, comp_feat_11_763, comp_feat_10_696, comp_feat_14_502, comp_feat_3_0, comp_feat_13_588, comp_feat_7_469, comp_feat_12_493, comp_feat_12_486, comp_feat_12_512, comp_feat_10_752, comp_feat_11_727, comp_feat_8_493, comp_feat_10_767, comp_feat_13_623, comp_feat_8_510, comp_feat_14_487, comp_feat_16_685, comp_feat_11_728, comp_feat_11_718, comp_feat_12_490, comp_feat_12_504, comp_feat_9_508, comp_feat_8_524, comp_feat_14_499, comp_feat_14_495, comp_feat_15_856, comp_feat_8_461, comp_feat_8_452, comp_feat_13_627, comp_feat_17_767, comp_feat_15_787, comp_feat_17_752, comp_feat_8_475, comp_feat_6_361, comp_feat_12_521, comp_feat_14_521, comp_feat_15_803, comp_feat_15_732, comp_feat_13_612, comp_feat_14_509, comp_feat_11_719, comp_feat_11_693, comp_feat_10_772, comp_feat_7_487, comp_feat_13_573, comp_feat_15_820, comp_feat_10_775, comp_feat_17_862, comp_feat_14_531, comp_feat_12_515, comp_feat_13_606, comp_feat_12_528, comp_feat_8_528, comp_feat_13_633, comp_feat_10_759, comp_feat_17_841, comp_feat_10_0, comp_feat_15_863, comp_feat_16_702, comp_feat_10_770, comp_feat_8_487, comp_feat_7_470, comp_feat_16_735, comp_feat_15_781, comp_feat_0_1, comp_feat_9_533, comp_feat_9_536, comp_feat_9_826, comp_feat_17_827, comp_feat_13_636, comp_feat_10_749, comp_feat_15_648, comp_feat_7_388, comp_feat_12_525, comp_feat_16_684, comp_feat_8_462, comp_feat_16_751, comp_feat_15_892, comp_feat_15_747, comp_feat_15_640, comp_feat_5_1, comp_feat_8_401, comp_feat_15_741, comp_feat_13_938, comp_feat_14_520, comp_feat_10_689, comp_feat_15_756, comp_feat_14_493, comp_feat_6_396, comp_feat_13_647, comp_feat_15_823, comp_feat_3_1, comp_feat_7_472, comp_feat_12_518, comp_feat_9_515, comp_feat_17_833, comp_feat_14_505, comp_feat_14_526, comp_feat_11_831, comp_feat_10_712, comp_feat_9_213, comp_feat_11_837, comp_feat_7_464, comp_feat_16_731, comp_feat_14_23, comp_feat_12_536, comp_feat_14_529, comp_feat_6_409, comp_feat_9_511, comp_feat_6_385, comp_feat_12_520, comp_feat_7_476, comp_feat_12_497, comp_feat_10_755, comp_feat_13_614, comp_feat_6_378, comp_feat_13_582, comp_feat_17_763, comp_feat_13_628, comp_feat_14_566, comp_feat_14_536, comp_feat_11_827, comp_feat_9_558, comp_feat_12_533, comp_feat_13_613, comp_feat_13_574, comp_feat_11_753, comp_feat_8_542, comp_feat_10_753, comp_feat_15_806, comp_feat_10_676, comp_feat_11_410, comp_feat_8_586, comp_feat_12_431, reg_decision
);


	assign reg_feat_8 = feat_8;

	assign reg_feat_13 = feat_13;

	assign reg_feat_10 = feat_10;

	assign reg_feat_12 = feat_12;

	assign reg_feat_2 = feat_2;

	assign reg_feat_14 = feat_14;

	assign reg_feat_9 = feat_9;

	assign reg_feat_11 = feat_11;

	assign reg_feat_17 = feat_17;

	assign reg_feat_16 = feat_16;

	assign reg_feat_5 = feat_5;

	assign reg_feat_0 = feat_0;

	assign reg_feat_1 = feat_1;

	assign reg_feat_6 = feat_6;

	assign reg_feat_7 = feat_7;

	assign reg_feat_3 = feat_3;

	assign reg_feat_15 = feat_15;

	assign decision = reg_decision;

endmodule


module COMPS(
KEY,
reg_feat_8, reg_feat_13, reg_feat_10, reg_feat_12, reg_feat_2, reg_feat_14, reg_feat_9, reg_feat_11, reg_feat_17, reg_feat_16, reg_feat_5, reg_feat_0, reg_feat_1, reg_feat_6, reg_feat_7, reg_feat_3, reg_feat_15, comp_feat_8_538, comp_feat_13_632, comp_feat_10_734, comp_feat_12_453, comp_feat_2_2, comp_feat_14_504, comp_feat_9_6, comp_feat_11_744, comp_feat_12_240, comp_feat_11_823, comp_feat_17_787, comp_feat_11_742, comp_feat_17_765, comp_feat_14_537, comp_feat_8_506, comp_feat_16_741, comp_feat_8_491, comp_feat_14_535, comp_feat_5_2, comp_feat_14_525, comp_feat_12_537, comp_feat_13_626, comp_feat_8_512, comp_feat_12_523, comp_feat_0_0, comp_feat_13_608, comp_feat_14_522, comp_feat_11_770, comp_feat_12_517, comp_feat_1_0, comp_feat_13_538, comp_feat_9_356, comp_feat_12_526, comp_feat_6_359, comp_feat_7_480, comp_feat_2_1, comp_feat_14_512, comp_feat_11_763, comp_feat_10_696, comp_feat_14_502, comp_feat_3_0, comp_feat_13_588, comp_feat_7_469, comp_feat_12_493, comp_feat_12_486, comp_feat_12_512, comp_feat_10_752, comp_feat_11_727, comp_feat_8_493, comp_feat_10_767, comp_feat_13_623, comp_feat_8_510, comp_feat_14_487, comp_feat_16_685, comp_feat_11_728, comp_feat_11_718, comp_feat_12_490, comp_feat_12_504, comp_feat_9_508, comp_feat_8_524, comp_feat_14_499, comp_feat_14_495, comp_feat_15_856, comp_feat_8_461, comp_feat_8_452, comp_feat_13_627, comp_feat_17_767, comp_feat_15_787, comp_feat_17_752, comp_feat_8_475, comp_feat_6_361, comp_feat_12_521, comp_feat_14_521, comp_feat_15_803, comp_feat_15_732, comp_feat_13_612, comp_feat_14_509, comp_feat_11_719, comp_feat_11_693, comp_feat_10_772, comp_feat_7_487, comp_feat_13_573, comp_feat_15_820, comp_feat_10_775, comp_feat_17_862, comp_feat_14_531, comp_feat_12_515, comp_feat_13_606, comp_feat_12_528, comp_feat_8_528, comp_feat_13_633, comp_feat_10_759, comp_feat_17_841, comp_feat_10_0, comp_feat_15_863, comp_feat_16_702, comp_feat_10_770, comp_feat_8_487, comp_feat_7_470, comp_feat_16_735, comp_feat_15_781, comp_feat_0_1, comp_feat_9_533, comp_feat_9_536, comp_feat_9_826, comp_feat_17_827, comp_feat_13_636, comp_feat_10_749, comp_feat_15_648, comp_feat_7_388, comp_feat_12_525, comp_feat_16_684, comp_feat_8_462, comp_feat_16_751, comp_feat_15_892, comp_feat_15_747, comp_feat_15_640, comp_feat_5_1, comp_feat_8_401, comp_feat_15_741, comp_feat_13_938, comp_feat_14_520, comp_feat_10_689, comp_feat_15_756, comp_feat_14_493, comp_feat_6_396, comp_feat_13_647, comp_feat_15_823, comp_feat_3_1, comp_feat_7_472, comp_feat_12_518, comp_feat_9_515, comp_feat_17_833, comp_feat_14_505, comp_feat_14_526, comp_feat_11_831, comp_feat_10_712, comp_feat_9_213, comp_feat_11_837, comp_feat_7_464, comp_feat_16_731, comp_feat_14_23, comp_feat_12_536, comp_feat_14_529, comp_feat_6_409, comp_feat_9_511, comp_feat_6_385, comp_feat_12_520, comp_feat_7_476, comp_feat_12_497, comp_feat_10_755, comp_feat_13_614, comp_feat_6_378, comp_feat_13_582, comp_feat_17_763, comp_feat_13_628, comp_feat_14_566, comp_feat_14_536, comp_feat_11_827, comp_feat_9_558, comp_feat_12_533, comp_feat_13_613, comp_feat_13_574, comp_feat_11_753, comp_feat_8_542, comp_feat_10_753, comp_feat_15_806, comp_feat_10_676, comp_feat_11_410, comp_feat_8_586, comp_feat_12_431
);
input [170:0] KEY;

input [9:0] reg_feat_8;
input [9:0] reg_feat_13;
input [9:0] reg_feat_10;
input [9:0] reg_feat_12;
input [1:0] reg_feat_2;
input [9:0] reg_feat_14;
input [9:0] reg_feat_9;
input [9:0] reg_feat_11;
input [9:0] reg_feat_17;
input [9:0] reg_feat_16;
input [1:0] reg_feat_5;
input [1:0] reg_feat_0;
input [0:0] reg_feat_1;
input [9:0] reg_feat_6;
input [9:0] reg_feat_7;
input [1:0] reg_feat_3;
input [9:0] reg_feat_15;
output [0:0] comp_feat_8_538;
output [0:0] comp_feat_13_632;
output [0:0] comp_feat_10_734;
output [0:0] comp_feat_12_453;
output [0:0] comp_feat_2_2;
output [0:0] comp_feat_14_504;
output [0:0] comp_feat_9_6;
output [0:0] comp_feat_11_744;
output [0:0] comp_feat_12_240;
output [0:0] comp_feat_11_823;
output [0:0] comp_feat_17_787;
output [0:0] comp_feat_11_742;
output [0:0] comp_feat_17_765;
output [0:0] comp_feat_14_537;
output [0:0] comp_feat_8_506;
output [0:0] comp_feat_16_741;
output [0:0] comp_feat_8_491;
output [0:0] comp_feat_14_535;
output [0:0] comp_feat_5_2;
output [0:0] comp_feat_14_525;
output [0:0] comp_feat_12_537;
output [0:0] comp_feat_13_626;
output [0:0] comp_feat_8_512;
output [0:0] comp_feat_12_523;
output [0:0] comp_feat_0_0;
output [0:0] comp_feat_13_608;
output [0:0] comp_feat_14_522;
output [0:0] comp_feat_11_770;
output [0:0] comp_feat_12_517;
output [0:0] comp_feat_1_0;
output [0:0] comp_feat_13_538;
output [0:0] comp_feat_9_356;
output [0:0] comp_feat_12_526;
output [0:0] comp_feat_6_359;
output [0:0] comp_feat_7_480;
output [0:0] comp_feat_2_1;
output [0:0] comp_feat_14_512;
output [0:0] comp_feat_11_763;
output [0:0] comp_feat_10_696;
output [0:0] comp_feat_14_502;
output [0:0] comp_feat_3_0;
output [0:0] comp_feat_13_588;
output [0:0] comp_feat_7_469;
output [0:0] comp_feat_12_493;
output [0:0] comp_feat_12_486;
output [0:0] comp_feat_12_512;
output [0:0] comp_feat_10_752;
output [0:0] comp_feat_11_727;
output [0:0] comp_feat_8_493;
output [0:0] comp_feat_10_767;
output [0:0] comp_feat_13_623;
output [0:0] comp_feat_8_510;
output [0:0] comp_feat_14_487;
output [0:0] comp_feat_16_685;
output [0:0] comp_feat_11_728;
output [0:0] comp_feat_11_718;
output [0:0] comp_feat_12_490;
output [0:0] comp_feat_12_504;
output [0:0] comp_feat_9_508;
output [0:0] comp_feat_8_524;
output [0:0] comp_feat_14_499;
output [0:0] comp_feat_14_495;
output [0:0] comp_feat_15_856;
output [0:0] comp_feat_8_461;
output [0:0] comp_feat_8_452;
output [0:0] comp_feat_13_627;
output [0:0] comp_feat_17_767;
output [0:0] comp_feat_15_787;
output [0:0] comp_feat_17_752;
output [0:0] comp_feat_8_475;
output [0:0] comp_feat_6_361;
output [0:0] comp_feat_12_521;
output [0:0] comp_feat_14_521;
output [0:0] comp_feat_15_803;
output [0:0] comp_feat_15_732;
output [0:0] comp_feat_13_612;
output [0:0] comp_feat_14_509;
output [0:0] comp_feat_11_719;
output [0:0] comp_feat_11_693;
output [0:0] comp_feat_10_772;
output [0:0] comp_feat_7_487;
output [0:0] comp_feat_13_573;
output [0:0] comp_feat_15_820;
output [0:0] comp_feat_10_775;
output [0:0] comp_feat_17_862;
output [0:0] comp_feat_14_531;
output [0:0] comp_feat_12_515;
output [0:0] comp_feat_13_606;
output [0:0] comp_feat_12_528;
output [0:0] comp_feat_8_528;
output [0:0] comp_feat_13_633;
output [0:0] comp_feat_10_759;
output [0:0] comp_feat_17_841;
output [0:0] comp_feat_10_0;
output [0:0] comp_feat_15_863;
output [0:0] comp_feat_16_702;
output [0:0] comp_feat_10_770;
output [0:0] comp_feat_8_487;
output [0:0] comp_feat_7_470;
output [0:0] comp_feat_16_735;
output [0:0] comp_feat_15_781;
output [0:0] comp_feat_0_1;
output [0:0] comp_feat_9_533;
output [0:0] comp_feat_9_536;
output [0:0] comp_feat_9_826;
output [0:0] comp_feat_17_827;
output [0:0] comp_feat_13_636;
output [0:0] comp_feat_10_749;
output [0:0] comp_feat_15_648;
output [0:0] comp_feat_7_388;
output [0:0] comp_feat_12_525;
output [0:0] comp_feat_16_684;
output [0:0] comp_feat_8_462;
output [0:0] comp_feat_16_751;
output [0:0] comp_feat_15_892;
output [0:0] comp_feat_15_747;
output [0:0] comp_feat_15_640;
output [0:0] comp_feat_5_1;
output [0:0] comp_feat_8_401;
output [0:0] comp_feat_15_741;
output [0:0] comp_feat_13_938;
output [0:0] comp_feat_14_520;
output [0:0] comp_feat_10_689;
output [0:0] comp_feat_15_756;
output [0:0] comp_feat_14_493;
output [0:0] comp_feat_6_396;
output [0:0] comp_feat_13_647;
output [0:0] comp_feat_15_823;
output [0:0] comp_feat_3_1;
output [0:0] comp_feat_7_472;
output [0:0] comp_feat_12_518;
output [0:0] comp_feat_9_515;
output [0:0] comp_feat_17_833;
output [0:0] comp_feat_14_505;
output [0:0] comp_feat_14_526;
output [0:0] comp_feat_11_831;
output [0:0] comp_feat_10_712;
output [0:0] comp_feat_9_213;
output [0:0] comp_feat_11_837;
output [0:0] comp_feat_7_464;
output [0:0] comp_feat_16_731;
output [0:0] comp_feat_14_23;
output [0:0] comp_feat_12_536;
output [0:0] comp_feat_14_529;
output [0:0] comp_feat_6_409;
output [0:0] comp_feat_9_511;
output [0:0] comp_feat_6_385;
output [0:0] comp_feat_12_520;
output [0:0] comp_feat_7_476;
output [0:0] comp_feat_12_497;
output [0:0] comp_feat_10_755;
output [0:0] comp_feat_13_614;
output [0:0] comp_feat_6_378;
output [0:0] comp_feat_13_582;
output [0:0] comp_feat_17_763;
output [0:0] comp_feat_13_628;
output [0:0] comp_feat_14_566;
output [0:0] comp_feat_14_536;
output [0:0] comp_feat_11_827;
output [0:0] comp_feat_9_558;
output [0:0] comp_feat_12_533;
output [0:0] comp_feat_13_613;
output [0:0] comp_feat_13_574;
output [0:0] comp_feat_11_753;
output [0:0] comp_feat_8_542;
output [0:0] comp_feat_10_753;
output [0:0] comp_feat_15_806;
output [0:0] comp_feat_10_676;
output [0:0] comp_feat_11_410;
output [0:0] comp_feat_8_586;
output [0:0] comp_feat_12_431;

wire [9:0] const_538_10;
assign const_538_10 = 10'b1000011010;
wire [9:0] const_632_10;
assign const_632_10 = 10'b1001111000;
wire [9:0] const_734_10;
assign const_734_10 = 10'b1011011110;
wire [9:0] const_453_10;
assign const_453_10 = 10'b0111000101;
wire [1:0] const_2_2;
assign const_2_2 = 2'b10;
wire [9:0] const_504_10;
assign const_504_10 = 10'b0111111000;
wire [9:0] const_6_10;
assign const_6_10 = 10'b0000000110;
wire [9:0] const_744_10;
assign const_744_10 = 10'b1011101000;
wire [9:0] const_240_10;
assign const_240_10 = 10'b0011110000;
wire [9:0] const_823_10;
assign const_823_10 = 10'b1100110111;
wire [9:0] const_787_10;
assign const_787_10 = 10'b1100010011;
wire [9:0] const_742_10;
assign const_742_10 = 10'b1011100110;
wire [9:0] const_765_10;
assign const_765_10 = 10'b1011111101;
wire [9:0] const_537_10;
assign const_537_10 = 10'b1000011001;
wire [9:0] const_506_10;
assign const_506_10 = 10'b0111111010;
wire [9:0] const_741_10;
assign const_741_10 = 10'b1011100101;
wire [9:0] const_491_10;
assign const_491_10 = 10'b0111101011;
wire [9:0] const_535_10;
assign const_535_10 = 10'b1000010111;
wire [9:0] const_525_10;
assign const_525_10 = 10'b1000001101;
wire [9:0] const_626_10;
assign const_626_10 = 10'b1001110010;
wire [9:0] const_512_10;
assign const_512_10 = 10'b1000000000;
wire [9:0] const_523_10;
assign const_523_10 = 10'b1000001011;
wire [1:0] const_0_2;
assign const_0_2 = 2'b00;
wire [9:0] const_608_10;
assign const_608_10 = 10'b1001100000;
wire [9:0] const_522_10;
assign const_522_10 = 10'b1000001010;
wire [9:0] const_770_10;
assign const_770_10 = 10'b1100000010;
wire [9:0] const_517_10;
assign const_517_10 = 10'b1000000101;
wire [0:0] const_0_1;
assign const_0_1 = 1'b0;
wire [9:0] const_356_10;
assign const_356_10 = 10'b0101100100;
wire [9:0] const_526_10;
assign const_526_10 = 10'b1000001110;
wire [9:0] const_359_10;
assign const_359_10 = 10'b0101100111;
wire [9:0] const_480_10;
assign const_480_10 = 10'b0111100000;
wire [1:0] const_1_2;
assign const_1_2 = 2'b01;
wire [9:0] const_763_10;
assign const_763_10 = 10'b1011111011;
wire [9:0] const_696_10;
assign const_696_10 = 10'b1010111000;
wire [9:0] const_502_10;
assign const_502_10 = 10'b0111110110;
wire [9:0] const_588_10;
assign const_588_10 = 10'b1001001100;
wire [9:0] const_469_10;
assign const_469_10 = 10'b0111010101;
wire [9:0] const_493_10;
assign const_493_10 = 10'b0111101101;
wire [9:0] const_486_10;
assign const_486_10 = 10'b0111100110;
wire [9:0] const_752_10;
assign const_752_10 = 10'b1011110000;
wire [9:0] const_727_10;
assign const_727_10 = 10'b1011010111;
wire [9:0] const_767_10;
assign const_767_10 = 10'b1011111111;
wire [9:0] const_623_10;
assign const_623_10 = 10'b1001101111;
wire [9:0] const_510_10;
assign const_510_10 = 10'b0111111110;
wire [9:0] const_487_10;
assign const_487_10 = 10'b0111100111;
wire [9:0] const_685_10;
assign const_685_10 = 10'b1010101101;
wire [9:0] const_728_10;
assign const_728_10 = 10'b1011011000;
wire [9:0] const_718_10;
assign const_718_10 = 10'b1011001110;
wire [9:0] const_490_10;
assign const_490_10 = 10'b0111101010;
wire [9:0] const_508_10;
assign const_508_10 = 10'b0111111100;
wire [9:0] const_524_10;
assign const_524_10 = 10'b1000001100;
wire [9:0] const_499_10;
assign const_499_10 = 10'b0111110011;
wire [9:0] const_495_10;
assign const_495_10 = 10'b0111101111;
wire [9:0] const_856_10;
assign const_856_10 = 10'b1101011000;
wire [9:0] const_461_10;
assign const_461_10 = 10'b0111001101;
wire [9:0] const_452_10;
assign const_452_10 = 10'b0111000100;
wire [9:0] const_627_10;
assign const_627_10 = 10'b1001110011;
wire [9:0] const_475_10;
assign const_475_10 = 10'b0111011011;
wire [9:0] const_361_10;
assign const_361_10 = 10'b0101101001;
wire [9:0] const_521_10;
assign const_521_10 = 10'b1000001001;
wire [9:0] const_803_10;
assign const_803_10 = 10'b1100100011;
wire [9:0] const_732_10;
assign const_732_10 = 10'b1011011100;
wire [9:0] const_612_10;
assign const_612_10 = 10'b1001100100;
wire [9:0] const_509_10;
assign const_509_10 = 10'b0111111101;
wire [9:0] const_719_10;
assign const_719_10 = 10'b1011001111;
wire [9:0] const_693_10;
assign const_693_10 = 10'b1010110101;
wire [9:0] const_772_10;
assign const_772_10 = 10'b1100000100;
wire [9:0] const_573_10;
assign const_573_10 = 10'b1000111101;
wire [9:0] const_820_10;
assign const_820_10 = 10'b1100110100;
wire [9:0] const_775_10;
assign const_775_10 = 10'b1100000111;
wire [9:0] const_862_10;
assign const_862_10 = 10'b1101011110;
wire [9:0] const_531_10;
assign const_531_10 = 10'b1000010011;
wire [9:0] const_515_10;
assign const_515_10 = 10'b1000000011;
wire [9:0] const_606_10;
assign const_606_10 = 10'b1001011110;
wire [9:0] const_528_10;
assign const_528_10 = 10'b1000010000;
wire [9:0] const_633_10;
assign const_633_10 = 10'b1001111001;
wire [9:0] const_759_10;
assign const_759_10 = 10'b1011110111;
wire [9:0] const_841_10;
assign const_841_10 = 10'b1101001001;
wire [9:0] const_0_10;
assign const_0_10 = 10'b0000000000;
wire [9:0] const_863_10;
assign const_863_10 = 10'b1101011111;
wire [9:0] const_702_10;
assign const_702_10 = 10'b1010111110;
wire [9:0] const_470_10;
assign const_470_10 = 10'b0111010110;
wire [9:0] const_735_10;
assign const_735_10 = 10'b1011011111;
wire [9:0] const_781_10;
assign const_781_10 = 10'b1100001101;
wire [9:0] const_533_10;
assign const_533_10 = 10'b1000010101;
wire [9:0] const_536_10;
assign const_536_10 = 10'b1000011000;
wire [9:0] const_826_10;
assign const_826_10 = 10'b1100111010;
wire [9:0] const_827_10;
assign const_827_10 = 10'b1100111011;
wire [9:0] const_636_10;
assign const_636_10 = 10'b1001111100;
wire [9:0] const_749_10;
assign const_749_10 = 10'b1011101101;
wire [9:0] const_648_10;
assign const_648_10 = 10'b1010001000;
wire [9:0] const_388_10;
assign const_388_10 = 10'b0110000100;
wire [9:0] const_684_10;
assign const_684_10 = 10'b1010101100;
wire [9:0] const_462_10;
assign const_462_10 = 10'b0111001110;
wire [9:0] const_751_10;
assign const_751_10 = 10'b1011101111;
wire [9:0] const_892_10;
assign const_892_10 = 10'b1101111100;
wire [9:0] const_747_10;
assign const_747_10 = 10'b1011101011;
wire [9:0] const_640_10;
assign const_640_10 = 10'b1010000000;
wire [9:0] const_401_10;
assign const_401_10 = 10'b0110010001;
wire [9:0] const_938_10;
assign const_938_10 = 10'b1110101010;
wire [9:0] const_520_10;
assign const_520_10 = 10'b1000001000;
wire [9:0] const_689_10;
assign const_689_10 = 10'b1010110001;
wire [9:0] const_756_10;
assign const_756_10 = 10'b1011110100;
wire [9:0] const_396_10;
assign const_396_10 = 10'b0110001100;
wire [9:0] const_647_10;
assign const_647_10 = 10'b1010000111;
wire [9:0] const_472_10;
assign const_472_10 = 10'b0111011000;
wire [9:0] const_518_10;
assign const_518_10 = 10'b1000000110;
wire [9:0] const_833_10;
assign const_833_10 = 10'b1101000001;
wire [9:0] const_505_10;
assign const_505_10 = 10'b0111111001;
wire [9:0] const_831_10;
assign const_831_10 = 10'b1100111111;
wire [9:0] const_712_10;
assign const_712_10 = 10'b1011001000;
wire [9:0] const_213_10;
assign const_213_10 = 10'b0011010101;
wire [9:0] const_837_10;
assign const_837_10 = 10'b1101000101;
wire [9:0] const_464_10;
assign const_464_10 = 10'b0111010000;
wire [9:0] const_731_10;
assign const_731_10 = 10'b1011011011;
wire [9:0] const_23_10;
assign const_23_10 = 10'b0000010111;
wire [9:0] const_529_10;
assign const_529_10 = 10'b1000010001;
wire [9:0] const_409_10;
assign const_409_10 = 10'b0110011001;
wire [9:0] const_511_10;
assign const_511_10 = 10'b0111111111;
wire [9:0] const_385_10;
assign const_385_10 = 10'b0110000001;
wire [9:0] const_476_10;
assign const_476_10 = 10'b0111011100;
wire [9:0] const_497_10;
assign const_497_10 = 10'b0111110001;
wire [9:0] const_755_10;
assign const_755_10 = 10'b1011110011;
wire [9:0] const_614_10;
assign const_614_10 = 10'b1001100110;
wire [9:0] const_378_10;
assign const_378_10 = 10'b0101111010;
wire [9:0] const_582_10;
assign const_582_10 = 10'b1001000110;
wire [9:0] const_628_10;
assign const_628_10 = 10'b1001110100;
wire [9:0] const_566_10;
assign const_566_10 = 10'b1000110110;
wire [9:0] const_558_10;
assign const_558_10 = 10'b1000101110;
wire [9:0] const_613_10;
assign const_613_10 = 10'b1001100101;
wire [9:0] const_574_10;
assign const_574_10 = 10'b1000111110;
wire [9:0] const_753_10;
assign const_753_10 = 10'b1011110001;
wire [9:0] const_542_10;
assign const_542_10 = 10'b1000011110;
wire [9:0] const_806_10;
assign const_806_10 = 10'b1100100110;
wire [9:0] const_676_10;
assign const_676_10 = 10'b1010100100;
wire [9:0] const_410_10;
assign const_410_10 = 10'b0110011010;
wire [9:0] const_586_10;
assign const_586_10 = 10'b1001001010;
wire [9:0] const_431_10;
assign const_431_10 = 10'b0110101111;

	assign comp_feat_8_538 = ((reg_feat_8 <= const_538_10)~^ KEY[0]);
	assign comp_feat_13_632 = (reg_feat_13 <= const_632_10);
	assign comp_feat_10_734 = (reg_feat_10 <= const_734_10);
	assign comp_feat_12_453 = ((reg_feat_12 <= const_453_10)~^ KEY[3]);
	assign comp_feat_2_2 = ((reg_feat_2 <= const_2_2)^ KEY[4]);
	assign comp_feat_14_504 = ((reg_feat_14 <= const_504_10)^ KEY[5]);
	assign comp_feat_9_6 = ((reg_feat_9 <= const_6_10)~^ KEY[6]);
	assign comp_feat_11_744 = ((reg_feat_11 <= const_744_10)^ KEY[7]);
	assign comp_feat_12_240 = ((reg_feat_12 <= const_240_10)~^ KEY[8]);
	assign comp_feat_11_823 = ((reg_feat_11 <= const_823_10)^ KEY[9]);
	assign comp_feat_17_787 = ((reg_feat_17 <= const_787_10)^ KEY[10]);
	assign comp_feat_11_742 = ((reg_feat_11 <= const_742_10)~^ KEY[11]);
	assign comp_feat_17_765 = ((reg_feat_17 <= const_765_10)^ KEY[12]);
	assign comp_feat_14_537 = (reg_feat_14 <= const_537_10);
	assign comp_feat_8_506 = ((reg_feat_8 <= const_506_10)^ KEY[14]);
	assign comp_feat_16_741 = ((reg_feat_16 <= const_741_10)~^ KEY[15]);
	assign comp_feat_8_491 = ((reg_feat_8 <= const_491_10)~^ KEY[16]);
	assign comp_feat_14_535 = ((reg_feat_14 <= const_535_10)~^ KEY[17]);
	assign comp_feat_5_2 = ((reg_feat_5 <= const_2_2)^ KEY[18]);
	assign comp_feat_14_525 = ((reg_feat_14 <= const_525_10)~^ KEY[19]);
	assign comp_feat_12_537 = ((reg_feat_12 <= const_537_10)^ KEY[20]);
	assign comp_feat_13_626 = ((reg_feat_13 <= const_626_10)^ KEY[21]);
	assign comp_feat_8_512 = ((reg_feat_8 <= const_512_10)~^ KEY[22]);
	assign comp_feat_12_523 = ((reg_feat_12 <= const_523_10)~^ KEY[23]);
	assign comp_feat_0_0 = ((reg_feat_0 <= const_0_2)~^ KEY[24]);
	assign comp_feat_13_608 = ((reg_feat_13 <= const_608_10)~^ KEY[25]);
	assign comp_feat_14_522 = (reg_feat_14 <= const_522_10);
	assign comp_feat_11_770 = (reg_feat_11 <= const_770_10);
	assign comp_feat_12_517 = (reg_feat_12 <= const_517_10);
	assign comp_feat_1_0 = ((reg_feat_1 <= const_0_1)^ KEY[29]);
	assign comp_feat_13_538 = ((reg_feat_13 <= const_538_10)^ KEY[30]);
	assign comp_feat_9_356 = ((reg_feat_9 <= const_356_10)^ KEY[31]);
	assign comp_feat_12_526 = ((reg_feat_12 <= const_526_10)~^ KEY[32]);
	assign comp_feat_6_359 = ((reg_feat_6 <= const_359_10)^ KEY[33]);
	assign comp_feat_7_480 = (reg_feat_7 <= const_480_10);
	assign comp_feat_2_1 = ((reg_feat_2 <= const_1_2)^ KEY[35]);
	assign comp_feat_14_512 = ((reg_feat_14 <= const_512_10)~^ KEY[36]);
	assign comp_feat_11_763 = (reg_feat_11 <= const_763_10);
	assign comp_feat_10_696 = ((reg_feat_10 <= const_696_10)~^ KEY[38]);
	assign comp_feat_14_502 = ((reg_feat_14 <= const_502_10)~^ KEY[39]);
	assign comp_feat_3_0 = ((reg_feat_3 <= const_0_2)~^ KEY[40]);
	assign comp_feat_13_588 = ((reg_feat_13 <= const_588_10)~^ KEY[41]);
	assign comp_feat_7_469 = (reg_feat_7 <= const_469_10);
	assign comp_feat_12_493 = ((reg_feat_12 <= const_493_10)~^ KEY[43]);
	assign comp_feat_12_486 = ((reg_feat_12 <= const_486_10)^ KEY[44]);
	assign comp_feat_12_512 = ((reg_feat_12 <= const_512_10)~^ KEY[45]);
	assign comp_feat_10_752 = ((reg_feat_10 <= const_752_10)^ KEY[46]);
	assign comp_feat_11_727 = ((reg_feat_11 <= const_727_10)^ KEY[47]);
	assign comp_feat_8_493 = ((reg_feat_8 <= const_493_10)~^ KEY[48]);
	assign comp_feat_10_767 = ((reg_feat_10 <= const_767_10)~^ KEY[49]);
	assign comp_feat_13_623 = (reg_feat_13 <= const_623_10);
	assign comp_feat_8_510 = ((reg_feat_8 <= const_510_10)~^ KEY[51]);
	assign comp_feat_14_487 = ((reg_feat_14 <= const_487_10)~^ KEY[52]);
	assign comp_feat_16_685 = ((reg_feat_16 <= const_685_10)~^ KEY[53]);
	assign comp_feat_11_728 = ((reg_feat_11 <= const_728_10)^ KEY[54]);
	assign comp_feat_11_718 = ((reg_feat_11 <= const_718_10)~^ KEY[55]);
	assign comp_feat_12_490 = ((reg_feat_12 <= const_490_10)~^ KEY[56]);
	assign comp_feat_12_504 = ((reg_feat_12 <= const_504_10)^ KEY[57]);
	assign comp_feat_9_508 = (reg_feat_9 <= const_508_10);
	assign comp_feat_8_524 = (reg_feat_8 <= const_524_10);
	assign comp_feat_14_499 = ((reg_feat_14 <= const_499_10)~^ KEY[60]);
	assign comp_feat_14_495 = ((reg_feat_14 <= const_495_10)^ KEY[61]);
	assign comp_feat_15_856 = ((reg_feat_15 <= const_856_10)^ KEY[62]);
	assign comp_feat_8_461 = ((reg_feat_8 <= const_461_10)^ KEY[63]);
	assign comp_feat_8_452 = ((reg_feat_8 <= const_452_10)^ KEY[64]);
	assign comp_feat_13_627 = ((reg_feat_13 <= const_627_10)^ KEY[65]);
	assign comp_feat_17_767 = ((reg_feat_17 <= const_767_10)^ KEY[66]);
	assign comp_feat_15_787 = ((reg_feat_15 <= const_787_10)^ KEY[67]);
	assign comp_feat_17_752 = ((reg_feat_17 <= const_752_10)~^ KEY[68]);
	assign comp_feat_8_475 = (reg_feat_8 <= const_475_10);
	assign comp_feat_6_361 = ((reg_feat_6 <= const_361_10)^ KEY[70]);
	assign comp_feat_12_521 = ((reg_feat_12 <= const_521_10)^ KEY[71]);
	assign comp_feat_14_521 = ((reg_feat_14 <= const_521_10)^ KEY[72]);
	assign comp_feat_15_803 = ((reg_feat_15 <= const_803_10)^ KEY[73]);
	assign comp_feat_15_732 = ((reg_feat_15 <= const_732_10)~^ KEY[74]);
	assign comp_feat_13_612 = ((reg_feat_13 <= const_612_10)~^ KEY[75]);
	assign comp_feat_14_509 = ((reg_feat_14 <= const_509_10)~^ KEY[76]);
	assign comp_feat_11_719 = (reg_feat_11 <= const_719_10);
	assign comp_feat_11_693 = ((reg_feat_11 <= const_693_10)^ KEY[78]);
	assign comp_feat_10_772 = ((reg_feat_10 <= const_772_10)~^ KEY[79]);
	assign comp_feat_7_487 = ((reg_feat_7 <= const_487_10)~^ KEY[80]);
	assign comp_feat_13_573 = ((reg_feat_13 <= const_573_10)^ KEY[81]);
	assign comp_feat_15_820 = ((reg_feat_15 <= const_820_10)~^ KEY[82]);
	assign comp_feat_10_775 = ((reg_feat_10 <= const_775_10)~^ KEY[83]);
	assign comp_feat_17_862 = ((reg_feat_17 <= const_862_10)~^ KEY[84]);
	assign comp_feat_14_531 = ((reg_feat_14 <= const_531_10)^ KEY[85]);
	assign comp_feat_12_515 = ((reg_feat_12 <= const_515_10)~^ KEY[86]);
	assign comp_feat_13_606 = (reg_feat_13 <= const_606_10);
	assign comp_feat_12_528 = ((reg_feat_12 <= const_528_10)~^ KEY[88]);
	assign comp_feat_8_528 = ((reg_feat_8 <= const_528_10)^ KEY[89]);
	assign comp_feat_13_633 = ((reg_feat_13 <= const_633_10)~^ KEY[90]);
	assign comp_feat_10_759 = ((reg_feat_10 <= const_759_10)^ KEY[91]);
	assign comp_feat_17_841 = ((reg_feat_17 <= const_841_10)~^ KEY[92]);
	assign comp_feat_10_0 = ((reg_feat_10 <= const_0_10)~^ KEY[93]);
	assign comp_feat_15_863 = ((reg_feat_15 <= const_863_10)~^ KEY[94]);
	assign comp_feat_16_702 = ((reg_feat_16 <= const_702_10)~^ KEY[95]);
	assign comp_feat_10_770 = ((reg_feat_10 <= const_770_10)~^ KEY[96]);
	assign comp_feat_8_487 = ((reg_feat_8 <= const_487_10)^ KEY[97]);
	assign comp_feat_7_470 = ((reg_feat_7 <= const_470_10)~^ KEY[98]);
	assign comp_feat_16_735 = ((reg_feat_16 <= const_735_10)~^ KEY[99]);
	assign comp_feat_15_781 = ((reg_feat_15 <= const_781_10)^ KEY[100]);
	assign comp_feat_0_1 = ((reg_feat_0 <= const_1_2)~^ KEY[101]);
	assign comp_feat_9_533 = ((reg_feat_9 <= const_533_10)~^ KEY[102]);
	assign comp_feat_9_536 = ((reg_feat_9 <= const_536_10)^ KEY[103]);
	assign comp_feat_9_826 = ((reg_feat_9 <= const_826_10)^ KEY[104]);
	assign comp_feat_17_827 = ((reg_feat_17 <= const_827_10)^ KEY[105]);
	assign comp_feat_13_636 = ((reg_feat_13 <= const_636_10)^ KEY[106]);
	assign comp_feat_10_749 = ((reg_feat_10 <= const_749_10)^ KEY[107]);
	assign comp_feat_15_648 = ((reg_feat_15 <= const_648_10)~^ KEY[108]);
	assign comp_feat_7_388 = ((reg_feat_7 <= const_388_10)~^ KEY[109]);
	assign comp_feat_12_525 = ((reg_feat_12 <= const_525_10)^ KEY[110]);
	assign comp_feat_16_684 = (reg_feat_16 <= const_684_10);
	assign comp_feat_8_462 = ((reg_feat_8 <= const_462_10)^ KEY[112]);
	assign comp_feat_16_751 = ((reg_feat_16 <= const_751_10)~^ KEY[113]);
	assign comp_feat_15_892 = ((reg_feat_15 <= const_892_10)~^ KEY[114]);
	assign comp_feat_15_747 = ((reg_feat_15 <= const_747_10)~^ KEY[115]);
	assign comp_feat_15_640 = ((reg_feat_15 <= const_640_10)~^ KEY[116]);
	assign comp_feat_5_1 = ((reg_feat_5 <= const_1_2)^ KEY[117]);
	assign comp_feat_8_401 = ((reg_feat_8 <= const_401_10)^ KEY[118]);
	assign comp_feat_15_741 = ((reg_feat_15 <= const_741_10)~^ KEY[119]);
	assign comp_feat_13_938 = (reg_feat_13 <= const_938_10);
	assign comp_feat_14_520 = ((reg_feat_14 <= const_520_10)~^ KEY[121]);
	assign comp_feat_10_689 = ((reg_feat_10 <= const_689_10)^ KEY[122]);
	assign comp_feat_15_756 = ((reg_feat_15 <= const_756_10)^ KEY[123]);
	assign comp_feat_14_493 = ((reg_feat_14 <= const_493_10)^ KEY[124]);
	assign comp_feat_6_396 = ((reg_feat_6 <= const_396_10)^ KEY[125]);
	assign comp_feat_13_647 = ((reg_feat_13 <= const_647_10)^ KEY[126]);
	assign comp_feat_15_823 = (reg_feat_15 <= const_823_10);
	assign comp_feat_3_1 = ((reg_feat_3 <= const_1_2)^ KEY[128]);
	assign comp_feat_7_472 = ((reg_feat_7 <= const_472_10)^ KEY[129]);
	assign comp_feat_12_518 = ((reg_feat_12 <= const_518_10)~^ KEY[130]);
	assign comp_feat_9_515 = ((reg_feat_9 <= const_515_10)^ KEY[131]);
	assign comp_feat_17_833 = ((reg_feat_17 <= const_833_10)~^ KEY[132]);
	assign comp_feat_14_505 = (reg_feat_14 <= const_505_10);
	assign comp_feat_14_526 = ((reg_feat_14 <= const_526_10)^ KEY[134]);
	assign comp_feat_11_831 = (reg_feat_11 <= const_831_10);
	assign comp_feat_10_712 = ((reg_feat_10 <= const_712_10)~^ KEY[136]);
	assign comp_feat_9_213 = (reg_feat_9 <= const_213_10);
	assign comp_feat_11_837 = ((reg_feat_11 <= const_837_10)~^ KEY[138]);
	assign comp_feat_7_464 = ((reg_feat_7 <= const_464_10)^ KEY[139]);
	assign comp_feat_16_731 = ((reg_feat_16 <= const_731_10)^ KEY[140]);
	assign comp_feat_14_23 = ((reg_feat_14 <= const_23_10)^ KEY[141]);
	assign comp_feat_12_536 = ((reg_feat_12 <= const_536_10)~^ KEY[142]);
	assign comp_feat_14_529 = ((reg_feat_14 <= const_529_10)^ KEY[143]);
	assign comp_feat_6_409 = (reg_feat_6 <= const_409_10);
	assign comp_feat_9_511 = ((reg_feat_9 <= const_511_10)~^ KEY[145]);
	assign comp_feat_6_385 = ((reg_feat_6 <= const_385_10)~^ KEY[146]);
	assign comp_feat_12_520 = ((reg_feat_12 <= const_520_10)~^ KEY[147]);
	assign comp_feat_7_476 = ((reg_feat_7 <= const_476_10)~^ KEY[148]);
	assign comp_feat_12_497 = ((reg_feat_12 <= const_497_10)^ KEY[149]);
	assign comp_feat_10_755 = (reg_feat_10 <= const_755_10);
	assign comp_feat_13_614 = ((reg_feat_13 <= const_614_10)~^ KEY[151]);
	assign comp_feat_6_378 = (reg_feat_6 <= const_378_10);
	assign comp_feat_13_582 = ((reg_feat_13 <= const_582_10)~^ KEY[153]);
	assign comp_feat_17_763 = ((reg_feat_17 <= const_763_10)^ KEY[154]);
	assign comp_feat_13_628 = ((reg_feat_13 <= const_628_10)^ KEY[155]);
	assign comp_feat_14_566 = ((reg_feat_14 <= const_566_10)^ KEY[156]);
	assign comp_feat_14_536 = (reg_feat_14 <= const_536_10);
	assign comp_feat_11_827 = ((reg_feat_11 <= const_827_10)^ KEY[158]);
	assign comp_feat_9_558 = ((reg_feat_9 <= const_558_10)~^ KEY[159]);
	assign comp_feat_12_533 = ((reg_feat_12 <= const_533_10)~^ KEY[160]);
	assign comp_feat_13_613 = ((reg_feat_13 <= const_613_10)^ KEY[161]);
	assign comp_feat_13_574 = ((reg_feat_13 <= const_574_10)^ KEY[162]);
	assign comp_feat_11_753 = ((reg_feat_11 <= const_753_10)^ KEY[163]);
	assign comp_feat_8_542 = ((reg_feat_8 <= const_542_10)^ KEY[164]);
	assign comp_feat_10_753 = ((reg_feat_10 <= const_753_10)^ KEY[165]);
	assign comp_feat_15_806 = ((reg_feat_15 <= const_806_10)^ KEY[166]);
	assign comp_feat_10_676 = (reg_feat_10 <= const_676_10);
	assign comp_feat_11_410 = ((reg_feat_11 <= const_410_10)~^ KEY[168]);
	assign comp_feat_8_586 = ((reg_feat_8 <= const_586_10)^ KEY[169]);
	assign comp_feat_12_431 = ((reg_feat_12 <= const_431_10)~^ KEY[170]);
endmodule


module ANDS(
comp_feat_8_538, comp_feat_13_632, comp_feat_10_734, comp_feat_12_453, comp_feat_2_2, comp_feat_14_504, comp_feat_9_6, comp_feat_11_744, comp_feat_12_240, comp_feat_11_823, comp_feat_17_787, comp_feat_11_742, comp_feat_17_765, comp_feat_14_537, comp_feat_8_506, comp_feat_16_741, comp_feat_8_491, comp_feat_14_535, comp_feat_5_2, comp_feat_14_525, comp_feat_12_537, comp_feat_13_626, comp_feat_8_512, comp_feat_12_523, comp_feat_0_0, comp_feat_13_608, comp_feat_14_522, comp_feat_11_770, comp_feat_12_517, comp_feat_1_0, comp_feat_13_538, comp_feat_9_356, comp_feat_12_526, comp_feat_6_359, comp_feat_7_480, comp_feat_2_1, comp_feat_14_512, comp_feat_11_763, comp_feat_10_696, comp_feat_14_502, comp_feat_3_0, comp_feat_13_588, comp_feat_7_469, comp_feat_12_493, comp_feat_12_486, comp_feat_12_512, comp_feat_10_752, comp_feat_11_727, comp_feat_8_493, comp_feat_10_767, comp_feat_13_623, comp_feat_8_510, comp_feat_14_487, comp_feat_16_685, comp_feat_11_728, comp_feat_11_718, comp_feat_12_490, comp_feat_12_504, comp_feat_9_508, comp_feat_8_524, comp_feat_14_499, comp_feat_14_495, comp_feat_15_856, comp_feat_8_461, comp_feat_8_452, comp_feat_13_627, comp_feat_17_767, comp_feat_15_787, comp_feat_17_752, comp_feat_8_475, comp_feat_6_361, comp_feat_12_521, comp_feat_14_521, comp_feat_15_803, comp_feat_15_732, comp_feat_13_612, comp_feat_14_509, comp_feat_11_719, comp_feat_11_693, comp_feat_10_772, comp_feat_7_487, comp_feat_13_573, comp_feat_15_820, comp_feat_10_775, comp_feat_17_862, comp_feat_14_531, comp_feat_12_515, comp_feat_13_606, comp_feat_12_528, comp_feat_8_528, comp_feat_13_633, comp_feat_10_759, comp_feat_17_841, comp_feat_10_0, comp_feat_15_863, comp_feat_16_702, comp_feat_10_770, comp_feat_8_487, comp_feat_7_470, comp_feat_16_735, comp_feat_15_781, comp_feat_0_1, comp_feat_9_533, comp_feat_9_536, comp_feat_9_826, comp_feat_17_827, comp_feat_13_636, comp_feat_10_749, comp_feat_15_648, comp_feat_7_388, comp_feat_12_525, comp_feat_16_684, comp_feat_8_462, comp_feat_16_751, comp_feat_15_892, comp_feat_15_747, comp_feat_15_640, comp_feat_5_1, comp_feat_8_401, comp_feat_15_741, comp_feat_13_938, comp_feat_14_520, comp_feat_10_689, comp_feat_15_756, comp_feat_14_493, comp_feat_6_396, comp_feat_13_647, comp_feat_15_823, comp_feat_3_1, comp_feat_7_472, comp_feat_12_518, comp_feat_9_515, comp_feat_17_833, comp_feat_14_505, comp_feat_14_526, comp_feat_11_831, comp_feat_10_712, comp_feat_9_213, comp_feat_11_837, comp_feat_7_464, comp_feat_16_731, comp_feat_14_23, comp_feat_12_536, comp_feat_14_529, comp_feat_6_409, comp_feat_9_511, comp_feat_6_385, comp_feat_12_520, comp_feat_7_476, comp_feat_12_497, comp_feat_10_755, comp_feat_13_614, comp_feat_6_378, comp_feat_13_582, comp_feat_17_763, comp_feat_13_628, comp_feat_14_566, comp_feat_14_536, comp_feat_11_827, comp_feat_9_558, comp_feat_12_533, comp_feat_13_613, comp_feat_13_574, comp_feat_11_753, comp_feat_8_542, comp_feat_10_753, comp_feat_15_806, comp_feat_10_676, comp_feat_11_410, comp_feat_8_586, comp_feat_12_431, reg_decision
);

input [0:0] comp_feat_8_538;
input [0:0] comp_feat_13_632;
input [0:0] comp_feat_10_734;
input [0:0] comp_feat_12_453;
input [0:0] comp_feat_2_2;
input [0:0] comp_feat_14_504;
input [0:0] comp_feat_9_6;
input [0:0] comp_feat_11_744;
input [0:0] comp_feat_12_240;
input [0:0] comp_feat_11_823;
input [0:0] comp_feat_17_787;
input [0:0] comp_feat_11_742;
input [0:0] comp_feat_17_765;
input [0:0] comp_feat_14_537;
input [0:0] comp_feat_8_506;
input [0:0] comp_feat_16_741;
input [0:0] comp_feat_8_491;
input [0:0] comp_feat_14_535;
input [0:0] comp_feat_5_2;
input [0:0] comp_feat_14_525;
input [0:0] comp_feat_12_537;
input [0:0] comp_feat_13_626;
input [0:0] comp_feat_8_512;
input [0:0] comp_feat_12_523;
input [0:0] comp_feat_0_0;
input [0:0] comp_feat_13_608;
input [0:0] comp_feat_14_522;
input [0:0] comp_feat_11_770;
input [0:0] comp_feat_12_517;
input [0:0] comp_feat_1_0;
input [0:0] comp_feat_13_538;
input [0:0] comp_feat_9_356;
input [0:0] comp_feat_12_526;
input [0:0] comp_feat_6_359;
input [0:0] comp_feat_7_480;
input [0:0] comp_feat_2_1;
input [0:0] comp_feat_14_512;
input [0:0] comp_feat_11_763;
input [0:0] comp_feat_10_696;
input [0:0] comp_feat_14_502;
input [0:0] comp_feat_3_0;
input [0:0] comp_feat_13_588;
input [0:0] comp_feat_7_469;
input [0:0] comp_feat_12_493;
input [0:0] comp_feat_12_486;
input [0:0] comp_feat_12_512;
input [0:0] comp_feat_10_752;
input [0:0] comp_feat_11_727;
input [0:0] comp_feat_8_493;
input [0:0] comp_feat_10_767;
input [0:0] comp_feat_13_623;
input [0:0] comp_feat_8_510;
input [0:0] comp_feat_14_487;
input [0:0] comp_feat_16_685;
input [0:0] comp_feat_11_728;
input [0:0] comp_feat_11_718;
input [0:0] comp_feat_12_490;
input [0:0] comp_feat_12_504;
input [0:0] comp_feat_9_508;
input [0:0] comp_feat_8_524;
input [0:0] comp_feat_14_499;
input [0:0] comp_feat_14_495;
input [0:0] comp_feat_15_856;
input [0:0] comp_feat_8_461;
input [0:0] comp_feat_8_452;
input [0:0] comp_feat_13_627;
input [0:0] comp_feat_17_767;
input [0:0] comp_feat_15_787;
input [0:0] comp_feat_17_752;
input [0:0] comp_feat_8_475;
input [0:0] comp_feat_6_361;
input [0:0] comp_feat_12_521;
input [0:0] comp_feat_14_521;
input [0:0] comp_feat_15_803;
input [0:0] comp_feat_15_732;
input [0:0] comp_feat_13_612;
input [0:0] comp_feat_14_509;
input [0:0] comp_feat_11_719;
input [0:0] comp_feat_11_693;
input [0:0] comp_feat_10_772;
input [0:0] comp_feat_7_487;
input [0:0] comp_feat_13_573;
input [0:0] comp_feat_15_820;
input [0:0] comp_feat_10_775;
input [0:0] comp_feat_17_862;
input [0:0] comp_feat_14_531;
input [0:0] comp_feat_12_515;
input [0:0] comp_feat_13_606;
input [0:0] comp_feat_12_528;
input [0:0] comp_feat_8_528;
input [0:0] comp_feat_13_633;
input [0:0] comp_feat_10_759;
input [0:0] comp_feat_17_841;
input [0:0] comp_feat_10_0;
input [0:0] comp_feat_15_863;
input [0:0] comp_feat_16_702;
input [0:0] comp_feat_10_770;
input [0:0] comp_feat_8_487;
input [0:0] comp_feat_7_470;
input [0:0] comp_feat_16_735;
input [0:0] comp_feat_15_781;
input [0:0] comp_feat_0_1;
input [0:0] comp_feat_9_533;
input [0:0] comp_feat_9_536;
input [0:0] comp_feat_9_826;
input [0:0] comp_feat_17_827;
input [0:0] comp_feat_13_636;
input [0:0] comp_feat_10_749;
input [0:0] comp_feat_15_648;
input [0:0] comp_feat_7_388;
input [0:0] comp_feat_12_525;
input [0:0] comp_feat_16_684;
input [0:0] comp_feat_8_462;
input [0:0] comp_feat_16_751;
input [0:0] comp_feat_15_892;
input [0:0] comp_feat_15_747;
input [0:0] comp_feat_15_640;
input [0:0] comp_feat_5_1;
input [0:0] comp_feat_8_401;
input [0:0] comp_feat_15_741;
input [0:0] comp_feat_13_938;
input [0:0] comp_feat_14_520;
input [0:0] comp_feat_10_689;
input [0:0] comp_feat_15_756;
input [0:0] comp_feat_14_493;
input [0:0] comp_feat_6_396;
input [0:0] comp_feat_13_647;
input [0:0] comp_feat_15_823;
input [0:0] comp_feat_3_1;
input [0:0] comp_feat_7_472;
input [0:0] comp_feat_12_518;
input [0:0] comp_feat_9_515;
input [0:0] comp_feat_17_833;
input [0:0] comp_feat_14_505;
input [0:0] comp_feat_14_526;
input [0:0] comp_feat_11_831;
input [0:0] comp_feat_10_712;
input [0:0] comp_feat_9_213;
input [0:0] comp_feat_11_837;
input [0:0] comp_feat_7_464;
input [0:0] comp_feat_16_731;
input [0:0] comp_feat_14_23;
input [0:0] comp_feat_12_536;
input [0:0] comp_feat_14_529;
input [0:0] comp_feat_6_409;
input [0:0] comp_feat_9_511;
input [0:0] comp_feat_6_385;
input [0:0] comp_feat_12_520;
input [0:0] comp_feat_7_476;
input [0:0] comp_feat_12_497;
input [0:0] comp_feat_10_755;
input [0:0] comp_feat_13_614;
input [0:0] comp_feat_6_378;
input [0:0] comp_feat_13_582;
input [0:0] comp_feat_17_763;
input [0:0] comp_feat_13_628;
input [0:0] comp_feat_14_566;
input [0:0] comp_feat_14_536;
input [0:0] comp_feat_11_827;
input [0:0] comp_feat_9_558;
input [0:0] comp_feat_12_533;
input [0:0] comp_feat_13_613;
input [0:0] comp_feat_13_574;
input [0:0] comp_feat_11_753;
input [0:0] comp_feat_8_542;
input [0:0] comp_feat_10_753;
input [0:0] comp_feat_15_806;
input [0:0] comp_feat_10_676;
input [0:0] comp_feat_11_410;
input [0:0] comp_feat_8_586;
input [0:0] comp_feat_12_431;
output [4:0] reg_decision;

wire [0:0] and_0;
wire [0:0] and_1;
wire [0:0] and_2;
wire [0:0] and_3;
wire [0:0] and_4;
wire [0:0] and_5;
wire [0:0] and_6;
wire [0:0] and_7;
wire [0:0] and_8;
wire [0:0] and_9;
wire [0:0] and_10;
wire [0:0] and_11;
wire [0:0] and_12;
wire [0:0] and_13;
wire [0:0] and_14;
wire [0:0] and_15;
wire [0:0] and_16;
wire [0:0] and_17;
wire [0:0] and_18;
wire [0:0] and_19;
wire [0:0] and_20;
wire [0:0] and_21;
wire [0:0] and_22;
wire [0:0] and_23;
wire [0:0] and_24;
wire [0:0] and_25;
wire [0:0] and_26;
wire [0:0] and_27;
wire [0:0] and_28;
wire [0:0] and_29;
wire [0:0] and_30;
wire [0:0] and_31;
wire [0:0] and_32;
wire [0:0] and_33;
wire [0:0] and_34;
wire [0:0] and_35;
wire [0:0] and_36;
wire [0:0] and_37;
wire [0:0] and_38;
wire [0:0] and_39;
wire [0:0] and_40;
wire [0:0] and_41;
wire [0:0] and_42;
wire [0:0] and_43;
wire [0:0] and_44;
wire [0:0] and_45;
wire [0:0] and_46;
wire [0:0] and_47;
wire [0:0] and_48;
wire [0:0] and_49;
wire [0:0] and_50;
wire [0:0] and_51;
wire [0:0] and_52;
wire [0:0] and_53;
wire [0:0] and_54;
wire [0:0] and_55;
wire [0:0] and_56;
wire [0:0] and_57;
wire [0:0] and_58;
wire [0:0] and_59;
wire [0:0] and_60;
wire [0:0] and_61;
wire [0:0] and_62;
wire [0:0] and_63;
wire [0:0] and_64;
wire [0:0] and_65;
wire [0:0] and_66;
wire [0:0] and_67;
wire [0:0] and_68;
wire [0:0] and_69;
wire [0:0] and_70;
wire [0:0] and_71;
wire [0:0] and_72;
wire [0:0] and_73;
wire [0:0] and_74;
wire [0:0] and_75;
wire [0:0] and_76;
wire [0:0] and_77;
wire [0:0] and_78;
wire [0:0] and_79;
wire [0:0] and_80;
wire [0:0] and_81;
wire [0:0] and_82;
wire [0:0] and_83;
wire [0:0] and_84;
wire [0:0] and_85;
wire [0:0] and_86;
wire [0:0] and_87;
wire [0:0] and_88;
wire [0:0] and_89;
wire [0:0] and_90;
wire [0:0] and_91;
wire [0:0] and_92;
wire [0:0] and_93;
wire [0:0] and_94;
wire [0:0] and_95;
wire [0:0] and_96;
wire [0:0] and_97;
wire [0:0] and_98;
wire [0:0] and_99;
wire [0:0] and_100;
wire [0:0] and_101;
wire [0:0] and_102;
wire [0:0] and_103;
wire [0:0] and_104;
wire [0:0] and_105;
wire [0:0] and_106;
wire [0:0] and_107;
wire [0:0] and_108;
wire [0:0] and_109;
wire [0:0] and_110;
wire [0:0] and_111;
wire [0:0] and_112;
wire [0:0] and_113;
wire [0:0] and_114;
wire [0:0] and_115;
wire [0:0] and_116;
wire [0:0] and_117;
wire [0:0] and_118;
wire [0:0] and_119;
wire [0:0] and_120;
wire [0:0] and_121;
wire [0:0] and_122;
wire [0:0] and_123;
wire [0:0] and_124;
wire [0:0] and_125;
wire [0:0] and_126;
wire [0:0] and_127;
wire [0:0] and_128;
wire [0:0] and_129;
wire [0:0] and_130;
wire [0:0] and_131;
wire [0:0] and_132;
wire [0:0] and_133;
wire [0:0] and_134;
wire [0:0] and_135;
wire [0:0] and_136;
wire [0:0] and_137;
wire [0:0] and_138;
wire [0:0] and_139;
wire [0:0] and_140;
wire [0:0] and_141;
wire [0:0] and_142;
wire [0:0] and_143;
wire [0:0] and_144;
wire [0:0] and_145;
wire [0:0] and_146;
wire [0:0] and_147;
wire [0:0] and_148;
wire [0:0] and_149;
wire [0:0] and_150;
wire [0:0] and_151;
wire [0:0] and_152;
wire [0:0] and_153;
wire [0:0] and_154;
wire [0:0] and_155;
wire [0:0] and_156;
wire [0:0] and_157;
wire [0:0] and_158;
wire [0:0] and_159;
wire [0:0] and_160;
wire [0:0] and_161;
wire [0:0] and_162;
wire [0:0] and_163;
wire [0:0] and_164;
wire [0:0] and_165;
wire [0:0] and_166;
wire [0:0] and_167;
wire [0:0] and_168;
wire [0:0] and_169;
wire [0:0] and_170;
wire [0:0] and_171;
wire [0:0] and_172;
wire [0:0] and_173;
wire [0:0] and_174;
wire [0:0] and_175;
wire [0:0] and_176;
wire [0:0] and_177;
wire [0:0] and_178;
wire [0:0] and_179;
wire [0:0] and_180;
wire [0:0] and_181;
wire [0:0] and_182;
wire [0:0] and_183;
wire [0:0] and_184;

assign and_0 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & comp_feat_14_525 & ~(comp_feat_12_537) & ~(comp_feat_8_512);

assign and_1 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & comp_feat_14_522 & ~(comp_feat_11_770) & comp_feat_1_0;

assign and_2 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & ~(comp_feat_14_522) & comp_feat_13_538 & ~(comp_feat_9_356);

assign and_3 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & ~(comp_feat_2_2) & ~(comp_feat_12_240);

assign and_4 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & ~(comp_feat_2_2) & ~(comp_feat_11_823);

assign and_5 = ~(comp_feat_8_538) & ~(comp_feat_16_735) & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & comp_feat_14_526 & comp_feat_11_831;

assign and_6 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & comp_feat_12_518 & ~(comp_feat_5_2);

assign and_7 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & ~(comp_feat_17_833);

assign and_8 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & comp_feat_14_505;

assign and_9 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & comp_feat_11_837 & comp_feat_7_464 & comp_feat_16_731 & ~(comp_feat_14_23);

assign and_10 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & comp_feat_11_837 & comp_feat_7_464 & ~(comp_feat_16_731) & ~(comp_feat_12_536);

assign and_11 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & comp_feat_11_837 & ~(comp_feat_7_464) & comp_feat_14_529 & ~(comp_feat_14_509);

assign and_12 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & comp_feat_11_837 & ~(comp_feat_7_464) & ~(comp_feat_14_529) & ~(comp_feat_6_409);

assign and_13 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & ~(comp_feat_11_837) & comp_feat_9_511;

assign and_14 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_9_515 & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & ~(comp_feat_13_614) & ~(comp_feat_6_378);

assign and_15 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_6_385 & comp_feat_12_520 & comp_feat_7_476 & comp_feat_12_497;

assign and_16 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_14_536 & ~(comp_feat_11_827);

assign and_17 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & ~(comp_feat_14_566) & ~(comp_feat_8_586);

assign reg_decision[0] = and_0 | and_1 | and_2 | and_3 | and_4 | and_5 | and_6 | and_7 | and_8 | and_9 | and_10 | and_11 | and_12 | and_13 | and_14 | and_15 | and_16 | and_17;

assign and_18 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & ~(comp_feat_14_525) & comp_feat_12_523 & comp_feat_0_0;

assign and_19 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & comp_feat_14_522 & ~(comp_feat_11_770) & ~(comp_feat_1_0);

assign and_20 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & ~(comp_feat_14_522) & comp_feat_13_538 & comp_feat_9_356;

assign and_21 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & comp_feat_12_526 & ~(comp_feat_6_359);

assign and_22 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & ~(comp_feat_12_526) & comp_feat_14_512 & ~(comp_feat_11_763);

assign and_23 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & comp_feat_2_2 & ~(comp_feat_14_504) & ~(comp_feat_11_744);

assign and_24 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_11_728) & ~(comp_feat_12_504) & ~(comp_feat_8_524);

assign and_25 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_14_499) & ~(comp_feat_8_461) & comp_feat_13_627;

assign and_26 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & comp_feat_7_469 & ~(comp_feat_12_493) & comp_feat_12_512;

assign and_27 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & comp_feat_10_767 & comp_feat_13_623 & comp_feat_8_510;

assign and_28 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & comp_feat_10_767 & ~(comp_feat_13_623) & ~(comp_feat_14_487);

assign and_29 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & ~(comp_feat_10_767) & comp_feat_16_685;

assign and_30 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & comp_feat_10_772 & ~(comp_feat_7_487) & ~(comp_feat_15_820);

assign and_31 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & ~(comp_feat_10_772) & ~(comp_feat_10_775) & ~(comp_feat_17_862);

assign and_32 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & comp_feat_7_487 & ~(comp_feat_14_531) & comp_feat_12_528;

assign and_33 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & ~(comp_feat_10_0) & comp_feat_15_863 & comp_feat_16_702 & comp_feat_8_461;

assign and_34 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & comp_feat_12_525 & comp_feat_16_684 & ~(comp_feat_8_462);

assign and_35 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & ~(comp_feat_15_640) & ~(comp_feat_8_401) & ~(comp_feat_13_938) & ~(comp_feat_14_520);

assign and_36 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_2_1 & ~(comp_feat_13_633) & ~(comp_feat_17_827) & comp_feat_10_689 & ~(comp_feat_15_756) & ~(comp_feat_14_493) & comp_feat_6_396;

assign and_37 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_2_1 & ~(comp_feat_13_633) & ~(comp_feat_17_827) & ~(comp_feat_10_689) & comp_feat_13_647 & ~(comp_feat_15_823);

assign and_38 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_2_1 & ~(comp_feat_13_633) & ~(comp_feat_17_827) & ~(comp_feat_10_689) & comp_feat_13_647 & comp_feat_3_1;

assign and_39 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & ~(comp_feat_17_841);

assign and_40 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_9_213) & comp_feat_11_837 & ~(comp_feat_7_464) & ~(comp_feat_14_529) & comp_feat_6_409;

assign and_41 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & ~(comp_feat_10_712) & ~(comp_feat_9_533);

assign and_42 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_9_515 & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & comp_feat_13_614;

assign and_43 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_6_385 & comp_feat_12_520 & comp_feat_7_476 & ~(comp_feat_12_497);

assign and_44 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_6_385 & ~(comp_feat_12_520) & ~(comp_feat_10_755) & comp_feat_13_628;

assign and_45 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_14_536 & comp_feat_11_827 & comp_feat_9_558 & comp_feat_12_533;

assign and_46 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_14_536) & comp_feat_13_613 & ~(comp_feat_13_574);

assign and_47 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_14_536) & ~(comp_feat_13_613) & ~(comp_feat_11_753);

assign and_48 = ~(comp_feat_8_538) & ~(comp_feat_12_537) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_10_753);

assign and_49 = ~(comp_feat_8_538) & ~(comp_feat_12_537) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_15_806 & ~(comp_feat_10_676);

assign and_50 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & ~(comp_feat_14_566) & comp_feat_8_586 & ~(comp_feat_12_431);

assign reg_decision[1] = and_18 | and_19 | and_20 | and_21 | and_22 | and_23 | and_24 | and_25 | and_26 | and_27 | and_28 | and_29 | and_30 | and_31 | and_32 | and_33 | and_34 | and_35 | and_36 | and_37 | and_38 | and_39 | and_40 | and_41 | and_42 | and_43 | and_44 | and_45 | and_46 | and_47 | and_48 | and_49 | and_50;

assign and_51 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & ~(comp_feat_17_765) & ~(comp_feat_8_491) & comp_feat_5_2;

assign and_52 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & ~(comp_feat_12_526) & ~(comp_feat_14_512) & ~(comp_feat_10_696);

assign and_53 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_8_506) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & ~(comp_feat_10_772) & comp_feat_10_775;

assign and_54 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_787 & comp_feat_17_752 & comp_feat_8_475;

assign and_55 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_787 & ~(comp_feat_17_752) & ~(comp_feat_6_361);

assign and_56 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_787) & comp_feat_12_521 & comp_feat_14_521;

assign and_57 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_787) & ~(comp_feat_12_521) & comp_feat_15_803;

assign and_58 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_732) & comp_feat_14_509 & ~(comp_feat_11_719);

assign and_59 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & comp_feat_2_2 & comp_feat_14_504 & comp_feat_9_6;

assign and_60 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_14_499 & comp_feat_14_495 & ~(comp_feat_15_856);

assign and_61 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_14_499) & comp_feat_8_461 & ~(comp_feat_8_452);

assign and_62 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & comp_feat_7_469 & comp_feat_12_493 & ~(comp_feat_12_486);

assign and_63 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & ~(comp_feat_7_469) & comp_feat_10_752 & ~(comp_feat_11_727);

assign and_64 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & ~(comp_feat_7_469) & ~(comp_feat_10_752) & ~(comp_feat_8_493);

assign and_65 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & comp_feat_10_767 & comp_feat_13_623 & ~(comp_feat_8_510);

assign and_66 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & comp_feat_10_772 & comp_feat_7_487 & ~(comp_feat_13_573);

assign and_67 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & comp_feat_14_531 & ~(comp_feat_12_515) & ~(comp_feat_13_606);

assign and_68 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & ~(comp_feat_14_531) & ~(comp_feat_12_528) & ~(comp_feat_8_528);

assign and_69 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & comp_feat_8_487 & ~(comp_feat_14_504) & comp_feat_7_470 & ~(comp_feat_16_735);

assign and_70 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & ~(comp_feat_8_487) & ~(comp_feat_15_781) & ~(comp_feat_0_1);

assign and_71 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & ~(comp_feat_10_770) & ~(comp_feat_9_533) & comp_feat_9_536;

assign and_72 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & ~(comp_feat_10_770) & ~(comp_feat_9_533) & ~(comp_feat_9_826);

assign and_73 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & ~(comp_feat_12_525) & comp_feat_16_751 & ~(comp_feat_15_892);

assign and_74 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & ~(comp_feat_12_525) & ~(comp_feat_16_751) & ~(comp_feat_15_747);

assign and_75 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_2_1 & ~(comp_feat_13_633) & ~(comp_feat_17_827) & ~(comp_feat_10_689) & comp_feat_13_647 & comp_feat_15_823 & ~(comp_feat_3_1);

assign and_76 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & ~(comp_feat_10_712) & comp_feat_9_533;

assign and_77 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_9_515) & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & ~(comp_feat_13_582) & ~(comp_feat_17_763);

assign and_78 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_14_536 & comp_feat_11_827 & comp_feat_9_558 & ~(comp_feat_12_533);

assign and_79 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_14_536) & ~(comp_feat_13_613) & comp_feat_11_753 & ~(comp_feat_8_542);

assign and_80 = ~(comp_feat_8_538) & ~(comp_feat_12_537) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_10_753 & ~(comp_feat_15_806);

assign reg_decision[2] = and_51 | and_52 | and_53 | and_54 | and_55 | and_56 | and_57 | and_58 | and_59 | and_60 | and_61 | and_62 | and_63 | and_64 | and_65 | and_66 | and_67 | and_68 | and_69 | and_70 | and_71 | and_72 | and_73 | and_74 | and_75 | and_76 | and_77 | and_78 | and_79 | and_80;

assign and_81 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & comp_feat_17_765 & ~(comp_feat_14_537) & comp_feat_16_741;

assign and_82 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & ~(comp_feat_17_765) & comp_feat_8_491 & ~(comp_feat_14_535);

assign and_83 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & comp_feat_14_525 & comp_feat_12_537 & comp_feat_13_626;

assign and_84 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & comp_feat_14_525 & ~(comp_feat_12_537) & comp_feat_8_512;

assign and_85 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & ~(comp_feat_14_525) & ~(comp_feat_12_523);

assign and_86 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & ~(comp_feat_14_525) & ~(comp_feat_0_0);

assign and_87 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & comp_feat_14_522 & comp_feat_11_770 & comp_feat_12_517;

assign and_88 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & ~(comp_feat_14_522) & ~(comp_feat_13_538);

assign and_89 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & comp_feat_12_526 & comp_feat_6_359 & comp_feat_7_480;

assign and_90 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & ~(comp_feat_12_526) & ~(comp_feat_14_512) & comp_feat_10_696;

assign and_91 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_787) & comp_feat_12_521 & ~(comp_feat_14_521);

assign and_92 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_787) & ~(comp_feat_12_521) & ~(comp_feat_15_803);

assign and_93 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & comp_feat_14_531 & comp_feat_12_515;

assign and_94 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_732 & comp_feat_13_612;

assign and_95 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & comp_feat_2_2 & comp_feat_14_504 & ~(comp_feat_9_6);

assign and_96 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & ~(comp_feat_2_2) & comp_feat_12_240 & comp_feat_11_823;

assign and_97 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_11_728 & ~(comp_feat_11_718) & comp_feat_12_490;

assign and_98 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_11_728) & comp_feat_12_504 & comp_feat_9_508;

assign and_99 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & comp_feat_7_469 & comp_feat_12_493 & comp_feat_12_486;

assign and_100 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & ~(comp_feat_7_469) & comp_feat_10_752 & comp_feat_11_727;

assign and_101 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & comp_feat_10_772 & comp_feat_7_487 & comp_feat_13_573;

assign and_102 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & comp_feat_14_531 & ~(comp_feat_12_515) & comp_feat_13_606;

assign and_103 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & ~(comp_feat_14_531) & ~(comp_feat_12_528) & comp_feat_8_528;

assign and_104 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & comp_feat_8_487 & ~(comp_feat_14_504) & comp_feat_7_470 & comp_feat_16_735;

assign and_105 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & comp_feat_10_749 & comp_feat_15_648;

assign and_106 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & comp_feat_10_749 & comp_feat_7_388;

assign and_107 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & comp_feat_12_525 & comp_feat_16_684 & comp_feat_8_462;

assign and_108 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & comp_feat_15_640 & comp_feat_5_1;

assign and_109 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & ~(comp_feat_15_640) & comp_feat_8_401 & comp_feat_15_741;

assign and_110 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_2_1 & ~(comp_feat_13_633) & ~(comp_feat_17_827) & comp_feat_10_689 & comp_feat_15_756;

assign and_111 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & comp_feat_17_841 & comp_feat_10_0;

assign and_112 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & comp_feat_17_841 & ~(comp_feat_15_863);

assign and_113 = ~(comp_feat_8_538) & comp_feat_16_735 & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & comp_feat_17_833 & ~(comp_feat_14_505);

assign and_114 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & comp_feat_12_518 & comp_feat_5_2 & comp_feat_9_515;

assign and_115 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & comp_feat_17_833 & ~(comp_feat_14_505) & ~(comp_feat_14_526);

assign and_116 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & ~(comp_feat_12_518) & comp_feat_17_833 & ~(comp_feat_14_505) & ~(comp_feat_11_831);

assign and_117 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & comp_feat_9_213;

assign and_118 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & comp_feat_11_837 & comp_feat_7_464 & comp_feat_16_731 & comp_feat_14_23;

assign and_119 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & comp_feat_11_837 & comp_feat_7_464 & ~(comp_feat_16_731) & comp_feat_12_536;

assign and_120 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & comp_feat_11_837 & ~(comp_feat_7_464) & comp_feat_14_529 & comp_feat_14_509;

assign and_121 = ~(comp_feat_8_538) & ~(comp_feat_15_781) & comp_feat_7_472 & comp_feat_10_712 & ~(comp_feat_11_837) & ~(comp_feat_9_511);

assign and_122 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_9_515) & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & comp_feat_13_582;

assign and_123 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_14_536) & comp_feat_13_613 & comp_feat_13_574;

assign and_124 = ~(comp_feat_8_538) & ~(comp_feat_12_537) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_10_753 & comp_feat_15_806 & comp_feat_10_676 & ~(comp_feat_11_410);

assign reg_decision[3] = and_81 | and_82 | and_83 | and_84 | and_85 | and_86 | and_87 | and_88 | and_89 | and_90 | and_91 | and_92 | and_93 | and_94 | and_95 | and_96 | and_97 | and_98 | and_99 | and_100 | and_101 | and_102 | and_103 | and_104 | and_105 | and_106 | and_107 | and_108 | and_109 | and_110 | and_111 | and_112 | and_113 | and_114 | and_115 | and_116 | and_117 | and_118 | and_119 | and_120 | and_121 | and_122 | and_123 | and_124;

assign and_125 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & comp_feat_17_765 & comp_feat_14_537;

assign and_126 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & comp_feat_17_765 & ~(comp_feat_16_741);

assign and_127 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & ~(comp_feat_17_765) & comp_feat_8_491 & comp_feat_14_535;

assign and_128 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & comp_feat_11_742 & ~(comp_feat_17_765) & ~(comp_feat_8_491) & ~(comp_feat_5_2);

assign and_129 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & comp_feat_17_787 & ~(comp_feat_11_742) & comp_feat_14_525 & comp_feat_12_537 & ~(comp_feat_13_626);

assign and_130 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & comp_feat_13_608 & comp_feat_14_522 & comp_feat_11_770 & ~(comp_feat_12_517);

assign and_131 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & comp_feat_12_526 & comp_feat_6_359 & ~(comp_feat_7_480);

assign and_132 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & ~(comp_feat_12_453) & ~(comp_feat_17_787) & ~(comp_feat_13_608) & ~(comp_feat_12_526) & comp_feat_14_512 & comp_feat_11_763;

assign and_133 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_8_506 & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & ~(comp_feat_10_772) & comp_feat_10_775;

assign and_134 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_787 & comp_feat_17_752 & ~(comp_feat_8_475);

assign and_135 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_5_2 & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_787 & ~(comp_feat_17_752) & comp_feat_6_361;

assign and_136 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & comp_feat_17_767 & comp_feat_15_732 & ~(comp_feat_13_612);

assign and_137 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_732) & ~(comp_feat_14_509);

assign and_138 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & comp_feat_17_767 & ~(comp_feat_15_732) & comp_feat_11_719;

assign and_139 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_5_2) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & comp_feat_14_531 & comp_feat_12_515;

assign and_140 = comp_feat_8_538 & comp_feat_13_632 & comp_feat_10_734 & comp_feat_12_453 & comp_feat_2_2 & ~(comp_feat_14_504) & comp_feat_11_744;

assign and_141 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_11_728 & comp_feat_11_718;

assign and_142 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_11_728 & ~(comp_feat_12_490);

assign and_143 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_11_728) & comp_feat_12_504 & ~(comp_feat_9_508);

assign and_144 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_13_626 & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_11_728) & ~(comp_feat_12_504) & comp_feat_8_524;

assign and_145 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_14_499 & ~(comp_feat_14_495);

assign and_146 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & comp_feat_14_499 & comp_feat_15_856;

assign and_147 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_14_499) & comp_feat_8_461 & comp_feat_8_452;

assign and_148 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_13_626) & comp_feat_14_502 & ~(comp_feat_3_0) & ~(comp_feat_14_499) & ~(comp_feat_8_461) & ~(comp_feat_13_627);

assign and_149 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & comp_feat_7_469 & ~(comp_feat_12_493) & ~(comp_feat_12_512);

assign and_150 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & comp_feat_13_588 & ~(comp_feat_7_469) & ~(comp_feat_10_752) & comp_feat_8_493;

assign and_151 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & comp_feat_10_767 & ~(comp_feat_13_623) & comp_feat_14_487;

assign and_152 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & comp_feat_14_502 & comp_feat_3_0 & ~(comp_feat_13_588) & ~(comp_feat_10_767) & ~(comp_feat_16_685);

assign and_153 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & comp_feat_10_772 & ~(comp_feat_7_487) & comp_feat_15_820;

assign and_154 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & comp_feat_11_693 & ~(comp_feat_10_772) & ~(comp_feat_10_775) & comp_feat_17_862;

assign and_155 = comp_feat_8_538 & comp_feat_13_632 & ~(comp_feat_10_734) & ~(comp_feat_14_502) & ~(comp_feat_17_767) & ~(comp_feat_11_693) & ~(comp_feat_7_487) & ~(comp_feat_14_531) & comp_feat_12_528;

assign and_156 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & comp_feat_17_841 & ~(comp_feat_10_0) & comp_feat_15_863 & ~(comp_feat_16_702);

assign and_157 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & comp_feat_10_759 & comp_feat_17_841 & ~(comp_feat_10_0) & comp_feat_15_863 & ~(comp_feat_8_461);

assign and_158 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & comp_feat_8_487 & comp_feat_14_504;

assign and_159 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & comp_feat_8_487 & ~(comp_feat_7_470);

assign and_160 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & ~(comp_feat_8_487) & comp_feat_15_781;

assign and_161 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & comp_feat_10_770 & ~(comp_feat_8_487) & comp_feat_0_1;

assign and_162 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & ~(comp_feat_10_770) & comp_feat_9_533;

assign and_163 = comp_feat_8_538 & ~(comp_feat_13_632) & comp_feat_13_633 & ~(comp_feat_10_759) & ~(comp_feat_10_770) & ~(comp_feat_9_536) & comp_feat_9_826;

assign and_164 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & comp_feat_10_749 & ~(comp_feat_15_648) & ~(comp_feat_7_388);

assign and_165 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & comp_feat_12_525 & ~(comp_feat_16_684);

assign and_166 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & ~(comp_feat_12_525) & comp_feat_16_751 & comp_feat_15_892;

assign and_167 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & comp_feat_13_636 & ~(comp_feat_10_749) & ~(comp_feat_12_525) & ~(comp_feat_16_751) & comp_feat_15_747;

assign and_168 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & comp_feat_15_640 & ~(comp_feat_5_1);

assign and_169 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & ~(comp_feat_15_640) & comp_feat_8_401 & ~(comp_feat_15_741);

assign and_170 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & ~(comp_feat_15_640) & ~(comp_feat_8_401) & comp_feat_13_938;

assign and_171 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & comp_feat_17_827 & ~(comp_feat_13_636) & ~(comp_feat_15_640) & ~(comp_feat_8_401) & comp_feat_14_520;

assign and_172 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & ~(comp_feat_17_827) & comp_feat_10_689 & ~(comp_feat_15_756) & comp_feat_14_493;

assign and_173 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & ~(comp_feat_17_827) & comp_feat_10_689 & ~(comp_feat_15_756) & ~(comp_feat_6_396);

assign and_174 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_13_633) & ~(comp_feat_17_827) & ~(comp_feat_10_689) & ~(comp_feat_13_647);

assign and_175 = comp_feat_8_538 & ~(comp_feat_13_632) & ~(comp_feat_2_1) & ~(comp_feat_13_633) & ~(comp_feat_17_827);

assign and_176 = ~(comp_feat_8_538) & comp_feat_15_781 & comp_feat_7_472 & comp_feat_12_518 & comp_feat_5_2 & ~(comp_feat_9_515);

assign and_177 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_9_515 & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & ~(comp_feat_13_614) & comp_feat_6_378;

assign and_178 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_9_515) & comp_feat_6_385 & ~(comp_feat_12_520) & comp_feat_10_755 & ~(comp_feat_13_582) & comp_feat_17_763;

assign and_179 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_6_385 & comp_feat_12_520 & ~(comp_feat_7_476);

assign and_180 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & comp_feat_6_385 & ~(comp_feat_12_520) & ~(comp_feat_10_755) & ~(comp_feat_13_628);

assign and_181 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_14_536 & comp_feat_11_827 & ~(comp_feat_9_558);

assign and_182 = ~(comp_feat_8_538) & comp_feat_12_537 & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & ~(comp_feat_14_536) & ~(comp_feat_13_613) & comp_feat_11_753 & comp_feat_8_542;

assign and_183 = ~(comp_feat_8_538) & ~(comp_feat_12_537) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & comp_feat_14_566 & comp_feat_10_753 & comp_feat_15_806 & comp_feat_10_676 & comp_feat_11_410;

assign and_184 = ~(comp_feat_8_538) & ~(comp_feat_7_472) & ~(comp_feat_6_385) & ~(comp_feat_14_566) & comp_feat_8_586 & comp_feat_12_431;

assign reg_decision[4] = and_125 | and_126 | and_127 | and_128 | and_129 | and_130 | and_131 | and_132 | and_133 | and_134 | and_135 | and_136 | and_137 | and_138 | and_139 | and_140 | and_141 | and_142 | and_143 | and_144 | and_145 | and_146 | and_147 | and_148 | and_149 | and_150 | and_151 | and_152 | and_153 | and_154 | and_155 | and_156 | and_157 | and_158 | and_159 | and_160 | and_161 | and_162 | and_163 | and_164 | and_165 | and_166 | and_167 | and_168 | and_169 | and_170 | and_171 | and_172 | and_173 | and_174 | and_175 | and_176 | and_177 | and_178 | and_179 | and_180 | and_181 | and_182 | and_183 | and_184;


endmodule
